module conversion(out_max, tens, ones);
 input[7:0] out_max;
 output[7:0] tens, ones;

 reg [7:0] tens, ones;

 
always @(out_max)
begin
case(out_max)
8'b00111111:   tens=8'h30;
8'b01000000:   tens=8'h30;
8'b01000001:   tens=8'h30;
8'b01000010:   tens=8'h30;
8'b01000011:   tens=8'h30;
8'b01000100:   tens=8'h30;
8'b01000101:   tens=8'h30;
8'b01000110:   tens=8'h30;
8'b01000111:   tens=8'h30;
8'b01001000:   tens=8'h30;
8'b01001001:   tens=8'h30;
8'b01001010:   tens=8'h30;
8'b01001011:   tens=8'h30;
8'b01001100:   tens=8'h30;
8'b01001101:   tens=8'h30;
8'b01001110:   tens=8'h30;
8'b01001111:   tens=8'h30;
8'b01010000:   tens=8'h30;
8'b01010001:   tens=8'h30;
8'b01010010:   tens=8'h30;
8'b01010011:   tens=8'h30;
8'b01010100:   tens=8'h30;
8'b01010101:   tens=8'h30;
8'b01010110:   tens=8'h30;
8'b01010111:   tens=8'h30;
8'b01011000:   tens=8'h30;
8'b01011001:   tens=8'h30;
8'b01011010:   tens=8'h30;
8'b01011011:   tens=8'h30;
8'b01011100:   tens=8'h30;
8'b01011101:   tens=8'h30;
8'b01011110:   tens=8'h30;
8'b01011111:   tens=8'h30;
8'b01100000:   tens=8'h30;
8'b01100001:   tens=8'h30;
8'b01100010:   tens=8'h30;
8'b01100011:   tens=8'h30;
8'b01100100:   tens=8'h30;
8'b01100101:   tens=8'h30;
8'b01100110:   tens=8'h30;
8'b01100111:   tens=8'h30;
8'b01101000:   tens=8'h30;
8'b01101001:   tens=8'h30;
8'b01101010:   tens=8'h30;
8'b01101011:   tens=8'h30;
8'b01101100:   tens=8'h30;
8'b01101101:   tens=8'h30;
8'b01101110:   tens=8'h30;
8'b01101111:   tens=8'h30;
8'b01110000:   tens=8'h30;
8'b01110001:   tens=8'h30;
8'b01110010:   tens=8'h30;
8'b01110011:   tens=8'h30;
8'b01110100:   tens=8'h30;
8'b01110101:   tens=8'h30;
8'b01110110:   tens=8'h30;
8'b01110111:   tens=8'h30;
8'b01111000:   tens=8'h30;
8'b01111001:   tens=8'h30;
8'b01111010:   tens=8'h30;
8'b01111011:   tens=8'h30;
8'b01111100:   tens=8'h30;
8'b01111101:   tens=8'h30;
8'b01111110:   tens=8'h30;
8'b01111111:   tens=8'h30;
8'b10000000:   tens=8'h30;
8'b10000001:   tens=8'h30;
8'b10000010:   tens=8'h30;
8'b10000011:   tens=8'h30;
8'b10000100:   tens=8'h30;
8'b10000101:   tens=8'h30;
8'b10000110:   tens=8'h30;
8'b10000111:   tens=8'h30;
8'b10001000:   tens=8'h30;
8'b10001001:   tens=8'h30;
8'b10001010:   tens=8'h30;
8'b10001011:   tens=8'h30;
8'b10001100:   tens=8'h30;
8'b10001101:   tens=8'h30;
8'b10001110:   tens=8'h30;
8'b10001111:   tens=8'h30;
8'b10010000:   tens=8'h30;
8'b10010001:   tens=8'h30;
8'b10010010:   tens=8'h30;
8'b10010011:   tens=8'h30;
8'b10010100:   tens=8'h30;
8'b10010101:   tens=8'h30;
8'b10010110:   tens=8'h30;
8'b10010111:   tens=8'h30;
8'b10011000:   tens=8'h30;
8'b10011001:   tens=8'h30;
8'b10011010:   tens=8'h30;
8'b10011011:   tens=8'h30;
8'b10011100:   tens=8'h30;
8'b10011101:   tens=8'h30;
8'b10011110:   tens=8'h30;
8'b10011111:   tens=8'h30;
8'b10100000:   tens=8'h30;
8'b10100001:   tens=8'h30;
8'b10100010:   tens=8'h30;
8'b10100011:   tens=8'h30;
8'b10100100:   tens=8'h30;
8'b10100101:   tens=8'h30;
8'b10100110:   tens=8'h30;
8'b10100111:   tens=8'h30;
8'b10101000:   tens=8'h30;
8'b10101001:   tens=8'h30;
8'b10101010:   tens=8'h30;
8'b10101011:   tens=8'h30;
8'b10101100:   tens=8'h30;
8'b10101101:   tens=8'h30;
8'b10101110:   tens=8'h30;
8'b10101111:   tens=8'h30;
8'b10110000:   tens=8'h30;
8'b10110001:   tens=8'h30;
8'b10110010:   tens=8'h30;
8'b10110011:   tens=8'h30;
8'b10110100:   tens=8'h30;
8'b10110101:   tens=8'h30;
8'b10110110:   tens=8'h30;
8'b10110110:   tens=8'h30;
8'b10110110:   tens=8'h30;
8'b10110110:   tens=8'h30;
8'b10111010:   tens=8'h30;
8'b10111011:   tens=8'h30;
8'b10111100:   tens=8'h30;
8'b10111101:   tens=8'h30;
8'b10111110:   tens=8'h31;
8'b10111111:   tens=8'h31;
8'b11000000:   tens=8'h31;
8'b11000001:   tens=8'h31;
8'b11000010:   tens=8'h31;
8'b11000011:   tens=8'h31;
8'b11000100:   tens=8'h31;
8'b11000101:   tens=8'h31;
8'b11000110:   tens=8'h31;
8'b11000111:   tens=8'h31;
8'b11001000:   tens=8'h31;
8'b11001001:   tens=8'h31;
8'b11001010:   tens=8'h31;
8'b11001011:   tens=8'h31;
8'b11001100:   tens=8'h31;
8'b11001101:   tens=8'h31;
8'b11001110:   tens=8'h31;
8'b11001111:   tens=8'h31;
8'b11010000:   tens=8'h31;
8'b11010001:   tens=8'h31;
8'b11010010:   tens=8'h31;
8'b11010011:   tens=8'h31;
8'b11010100:   tens=8'h31;
8'b11010101:   tens=8'h31;
8'b11010110:   tens=8'h31;
8'b11010111:   tens=8'h31;
8'b11011000:   tens=8'h31;
8'b11011001:   tens=8'h31;
8'b11011010:   tens=8'h31;
8'b11011011:   tens=8'h31;
8'b	11011101	:	tens=	8'h	31	;
8'b	11011110	:	tens=	8'h	31	;
8'b	11011111	:	tens=	8'h	32	;
8'b	11100000	:	tens=	8'h	32	;
8'b	11100001	:	tens=	8'h	32	;
8'b	11100010	:	tens=	8'h	32	;
8'b	11100011	:	tens=	8'h	32	;
8'b	11100100	:	tens=	8'h	32	;
8'b	11100101	:	tens=	8'h	32	;
8'b	11100110	:	tens=	8'h	33	;
8'b	11100111	:	tens=	8'h	33	;
8'b	11101000	:	tens=	8'h	33	;
8'b	11101001	:	tens=	8'h	33	;
8'b	11101010	:	tens=	8'h	33	;
8'b	11101011	:	tens=	8'h	34	;
8'b	11101100	:	tens=	8'h	34	;
8'b	11101101	:	tens=	8'h	34	;
8'b	11101110	:	tens=	8'h	35	;
8'b	11101111	:	tens=	8'h	36	;
8'b	11110000	:	tens=	8'h	38	;
8'b	11110001	:	tens=	8'h	38	;
8'b	11110010	:	tens=	8'h	38	;
8'b	11110011	:	tens=	8'h	38	;
8'b	11110100	:	tens=	8'h	38	;
8'b	11110101	:	tens=	8'h	38	;
8'b	11110110	:	tens=	8'h	38	;
8'b	11110111	:	tens=	8'h	38	;
8'b	11111000	:	tens=	8'h	38	;
8'b	11111001	:	tens=	8'h	39	;
8'b	11111010	:	tens=	8'h	39	;
8'b	11111011	:	tens=	8'h	39	;
8'b	11111100	:	tens=	8'h	39	;
8'b	11111101	:	tens=	8'h	39	;
8'b	11111110	:	tens=	8'h	39	;
8'b	11111111	:	tens=	8'h	39	;

default: tens=8'h30;
endcase

case(out_max)
8'b00111111:   ones=8'h31;
8'b01000000:   ones=8'h31;
8'b01000001:   ones=8'h31;
8'b01000010:   ones=8'h31;
8'b01000011:   ones=8'h31;
8'b01000100:   ones=8'h31;
8'b01000101:   ones=8'h31;
8'b01000110:   ones=8'h31;
8'b01000111:   ones=8'h31;
8'b01001000:   ones=8'h31;
8'b01001001:   ones=8'h31;
8'b01001010:   ones=8'h31;
8'b01001011:   ones=8'h31;
8'b01001100:   ones=8'h31;
8'b01001101:   ones=8'h31;
8'b01001110:   ones=8'h31;
8'b01001111:   ones=8'h31;
8'b01010000:   ones=8'h31;
8'b01010001:   ones=8'h31;
8'b01010010:   ones=8'h31;
8'b01010011:   ones=8'h31;
8'b01010100:   ones=8'h31;
8'b01010101:   ones=8'h31;
8'b01010110:   ones=8'h31;
8'b01010111:   ones=8'h31;
8'b01011000:   ones=8'h31;
8'b01011001:   ones=8'h31;
8'b01011010:   ones=8'h31;
8'b01011011:   ones=8'h31;
8'b01011100:   ones=8'h31;
8'b01011101:   ones=8'h31;
8'b01011110:   ones=8'h31;
8'b01011111:   ones=8'h31;
8'b01100000:   ones=8'h31;
8'b01100001:   ones=8'h31;
8'b01100010:   ones=8'h31;
8'b01100011:   ones=8'h31;
8'b01100100:   ones=8'h31;
8'b01100101:   ones=8'h31;
8'b01100110:   ones=8'h31;
8'b01100111:   ones=8'h31;
8'b01101000:   ones=8'h31;
8'b01101001:   ones=8'h31;
8'b01101010:   ones=8'h31;
8'b01101011:   ones=8'h32;
8'b01101100:   ones=8'h32;
8'b01101101:   ones=8'h32;
8'b01101110:   ones=8'h32;
8'b01101111:   ones=8'h32;
8'b01110000:   ones=8'h32;
8'b01110001:   ones=8'h32;
8'b01110010:   ones=8'h32;
8'b01110011:   ones=8'h32;
8'b01110100:   ones=8'h32;
8'b01110101:   ones=8'h32;
8'b01110110:   ones=8'h32;
8'b01110111:   ones=8'h32;
8'b01111000:   ones=8'h32;
8'b01111001:   ones=8'h32;
8'b01111010:   ones=8'h32;
8'b01111011:   ones=8'h32;
8'b01111100:   ones=8'h32;
8'b01111101:   ones=8'h33;
8'b01111110:   ones=8'h33;
8'b01111111:   ones=8'h33;
8'b10000000:   ones=8'h33;
8'b10000001:   ones=8'h33;
8'b10000010:   ones=8'h33;
8'b10000011:   ones=8'h33;
8'b10000100:   ones=8'h33;
8'b10000101:   ones=8'h33;
8'b10000110:   ones=8'h33;
8'b10000111:   ones=8'h33;
8'b10001000:   ones=8'h34;
8'b10001001:   ones=8'h34;
8'b10001010:   ones=8'h34;
8'b10001011:   ones=8'h34;
8'b10001100:   ones=8'h34;
8'b10001101:   ones=8'h34;
8'b10001110:   ones=8'h34;
8'b10001111:   ones=8'h34;
8'b10010000:   ones=8'h34;
8'b10010001:   ones=8'h34;
8'b10010010:   ones=8'h34;
8'b10010011:   ones=8'h34;
8'b10010100:   ones=8'h34;
8'b10010101:   ones=8'h34;
8'b10010110:   ones=8'h34;
8'b10010111:   ones=8'h34;
8'b10011000:   ones=8'h35;
8'b10011001:   ones=8'h35;
8'b10011010:   ones=8'h35;
8'b10011011:   ones=8'h35;
8'b10011100:   ones=8'h35;
8'b10011101:   ones=8'h35;
8'b10011110:   ones=8'h35;
8'b10011111:   ones=8'h35;
8'b10100000:   ones=8'h35;
8'b10100001:   ones=8'h35;
8'b10100010:   ones=8'h35;
8'b10100011:   ones=8'h35;
8'b10100100:   ones=8'h35;
8'b10100101:   ones=8'h36;
8'b10100110:   ones=8'h36;
8'b10100111:   ones=8'h36;
8'b10101000:   ones=8'h36;
8'b10101001:   ones=8'h36;
8'b10101010:   ones=8'h36;
8'b10101011:   ones=8'h36;
8'b10101100:   ones=8'h36;
8'b10101101:   ones=8'h36;
8'b10101110:   ones=8'h36;
8'b10101111:   ones=8'h36;
8'b10110000:   ones=8'h36;
8'b10110001:   ones=8'h36;
8'b10110010:   ones=8'h36;
8'b10110011:   ones=8'h36;
8'b10110100:   ones=8'h37;
8'b10110101:   ones=8'h37;
8'b10110110:   ones=8'h38;
8'b10110110:   ones=8'h38;
8'b10110110:   ones=8'h38;
8'b10110110:   ones=8'h39;
8'b10111010:   ones=8'h39;
8'b10111011:   ones=8'h39;
8'b10111100:   ones=8'h39;
8'b10111101:   ones=8'h39;
8'b	10111110	:	ones=	8'h	30	;
8'b	10111111	:	ones=	8'h	30	;
8'b	11000000	:	ones=	8'h	30	;
8'b	11000001	:	ones=	8'h	30	;
8'b	11000010	:	ones=	8'h	30	;
8'b	11000011	:	ones=	8'h	31	;
8'b	11000100	:	ones=	8'h	31	;
8'b	11000101	:	ones=	8'h	31	;
8'b	11000110	:	ones=	8'h	31	;
8'b	11000111	:	ones=	8'h	31	;
8'b	11001000	:	ones=	8'h	32	;
8'b	11001001	:	ones=	8'h	32	;
8'b	11001010	:	ones=	8'h	32	;
8'b	11001011	:	ones=	8'h	32	;
8'b	11001100	:	ones=	8'h	32	;
8'b	11001101	:	ones=	8'h	33	;
8'b	11001110	:	ones=	8'h	33	;
8'b	11001111	:	ones=	8'h	33	;
8'b	11010000	:	ones=	8'h	33	;
8'b	11010001	:	ones=	8'h	33	;
8'b	11010010	:	ones=	8'h	34	;
8'b	11010011	:	ones=	8'h	34	;
8'b	11010100	:	ones=	8'h	34	;
8'b	11010101	:	ones=	8'h	34	;
8'b	11010110	:	ones=	8'h	34	;
8'b	11010111	:	ones=	8'h	34	;
8'b	11011000	:	ones=	8'h	34	;
8'b	11011001	:	ones=	8'h	34	;
8'b	11011010	:	ones=	8'h	34	;
8'b	11011011	:	ones=	8'h	34	;
8'b	11011100	:	ones=	8'h	35	;
8'b	11011101	:	ones=	8'h	37	;
8'b	11011110	:	ones=	8'h	38	;
8'b	11011111	:	ones=	8'h	30	;
8'b	11100000	:	ones=	8'h	31	;
8'b	11100001	:	ones=	8'h	33	;
8'b	11100010	:	ones=	8'h	35	;
8'b	11100011	:	ones=	8'h	36	;
8'b	11100100	:	ones=	8'h	38	;
8'b	11100101	:	ones=	8'h	39	;
8'b	11100110	:	ones=	8'h	31	;
8'b	11100111	:	ones=	8'h	33	;
8'b	11101000	:	ones=	8'h	34	;
8'b	11101001	:	ones=	8'h	36	;
8'b	11101010	:	ones=	8'h	38	;
8'b	11101011	:	ones=	8'h	31	;
8'b	11101100	:	ones=	8'h	34	;
8'b	11101101	:	ones=	8'h	38	;
8'b	11101110	:	ones=	8'h	37	;
8'b	11101111	:	ones=	8'h	38	;
8'b	11110000	:	ones=	8'h	31	;
8'b	11110001	:	ones=	8'h	32	;
8'b	11110010	:	ones=	8'h	33	;
8'b	11110011	:	ones=	8'h	34	;
8'b	11110100	:	ones=	8'h	35	;
8'b	11110101	:	ones=	8'h	36	;
8'b	11110110	:	ones=	8'h	37	;
8'b	11110111	:	ones=	8'h	38	;
8'b	11111000	:	ones=	8'h	39	;
8'b	11111001	:	ones=	8'h	30	;
8'b	11111010	:	ones=	8'h	31	;
8'b	11111011	:	ones=	8'h	32	;

default: ones=8'h30;
endcase
end

endmodule